module	sprite_storage	(	
//		--------	Clock Input	 	
					input		logic	clk,
					input		logic	resetN,
					input    logic frame_start,
					input    logic [0:10] requested_x,
					input    logic [0:10] requested_y,
					input    logic [0:7] ai_car_color,
					input    logic [0:7] player_car_color,
					input    logic [0:7] bg_color,
					input    logic [0:7] fl_color,
					output	logic [0:16*16-1][7:0] out_car1,
					output	logic [0:16*16-1][7:0] out_car2,
					output	logic [0:16*16-1][7:0] out_car3,
					output	logic [0:16*16-1][7:0] out_ai_car_red,
					output	logic [0:16*16-1][7:0] out_ai_car_yellow,
					output	logic [0:32*128-1][7:0] out_background,
					output	logic [0:16*16-1][7:0] out_finish_line,
					output	logic	[7:0] RGBout,  //rgb value from the bitmap 
					output   logic [0:1] collisions
);

const logic[0:15][0:15][7:0] car1 = {
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'he4,8'he4,8'h00,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'he4,8'he4,8'he4,8'hc0,8'h00,8'h62,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'he4,8'he4,8'he4,8'hc0,8'hc0,8'h62,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'he4,8'hff,8'he4,8'he4,8'he4,8'he4,8'hc0,8'hc0,8'h00,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'he4,8'hff,8'he4,8'he4,8'h00,8'he4,8'hc0,8'hc0,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'he4,8'hff,8'he4,8'h00,8'h00,8'h00,8'hc0,8'hc0,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'he4,8'he4,8'h00,8'h00,8'h00,8'h00,8'hc0,8'hc0,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'h00,8'he4,8'he4,8'he4,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'h00,8'hff,8'he4,8'he4,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'h00,8'hff,8'he4,8'he4,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'h00,8'h00,8'h00,8'h00,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'he4,8'he4,8'hff,8'h00,8'h00,8'h00,8'hc0,8'hc0,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'he4,8'h00,8'he4,8'he4,8'he4,8'he4,8'h00,8'hc0,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'he4,8'h00,8'he4,8'he4,8'he4,8'he4,8'h00,8'hc0,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hc0,8'hc0,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'he4,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hc0,8'h00,8'h62,8'h62,8'h62}};

const logic[0:15][0:15][7:0] car2 = {
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'he4,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'hff,8'he4,8'he4,8'he4,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'he4,8'hff,8'he4,8'he4,8'he4,8'he4,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'hff,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'he4,8'h00,8'h00,8'he4,8'he4,8'he4,8'he4,8'he4,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'he4,8'hff,8'h00,8'h00,8'h00,8'he4,8'he4,8'he4,8'he4,8'h62},
	{8'h62,8'h62,8'h62,8'he4,8'hff,8'he4,8'hff,8'he4,8'he4,8'h00,8'h00,8'h00,8'he4,8'he4,8'h00,8'h62},
	{8'h62,8'h62,8'he4,8'hff,8'he4,8'h00,8'h00,8'he4,8'he4,8'he4,8'h00,8'he4,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'he4,8'he4,8'he4,8'he4,8'h00,8'h00,8'h00,8'he4,8'hc0,8'hc0,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'he4,8'he4,8'he4,8'he4,8'he4,8'h00,8'h00,8'hc0,8'hc0,8'h00,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h00,8'h00,8'he4,8'he4,8'he4,8'he4,8'h00,8'hc0,8'hc0,8'hc0,8'h00,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h00,8'he4,8'he4,8'he4,8'he4,8'hc0,8'hc0,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h00,8'he4,8'he4,8'he4,8'hc0,8'hc0,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h00,8'he4,8'he4,8'he4,8'hc0,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h00,8'he4,8'he4,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'h00,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62}};

const logic[0:15][0:15][7:0] car3 = {
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'he4,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'he4,8'hff,8'hff,8'he4,8'he4,8'he4,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'h62,8'he4,8'hff,8'he4,8'he4,8'he4,8'he4,8'he4,8'h62},
	{8'h62,8'h62,8'h62,8'he4,8'he4,8'he4,8'hff,8'he4,8'he4,8'h00,8'he4,8'he4,8'he4,8'he4,8'he4,8'h62},
	{8'h62,8'h62,8'he4,8'he4,8'hff,8'he4,8'he4,8'he4,8'h00,8'h00,8'h00,8'he4,8'he4,8'he4,8'he4,8'h62},
	{8'h62,8'he4,8'he4,8'hff,8'h00,8'h00,8'he4,8'he4,8'he4,8'h00,8'h00,8'he4,8'he4,8'he4,8'he4,8'h62},
	{8'h00,8'he4,8'he4,8'he4,8'he4,8'h00,8'h00,8'he4,8'he4,8'h00,8'h00,8'he4,8'he4,8'hc0,8'h00,8'h62},
	{8'h00,8'he4,8'he4,8'he4,8'he4,8'h00,8'h00,8'h00,8'he4,8'he4,8'he4,8'hc0,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h00,8'h00,8'he4,8'he4,8'he4,8'h00,8'h00,8'he4,8'hc0,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h00,8'he4,8'he4,8'he4,8'h00,8'h00,8'he4,8'hc0,8'h00,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h00,8'he4,8'he4,8'he4,8'he4,8'he4,8'h00,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h00,8'he4,8'he4,8'he4,8'he4,8'hc0,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h00,8'he4,8'he4,8'he4,8'hc0,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h00,8'he4,8'he4,8'h00,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62}};

	
const logic[0:15][0:15][7:0] ai_car_red = {
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'he4,8'hff,8'he4,8'he4,8'he4,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'hff,8'he4,8'he4,8'he4,8'he4,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'hff,8'he4,8'he4,8'he4,8'he4,8'he4,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'hff,8'he4,8'he4,8'he4,8'he4,8'he4,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'hff,8'he4,8'he4,8'he4,8'he4,8'he4,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'hff,8'h00,8'h00,8'h00,8'he4,8'he4,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'h91,8'h00,8'h00,8'h00,8'h00,8'he4,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'h00,8'he4,8'he4,8'he4,8'h00,8'he4,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'h00,8'he4,8'he4,8'he4,8'h00,8'he4,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'h00,8'he4,8'he4,8'he4,8'h00,8'he4,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'h00,8'he4,8'he4,8'he4,8'h00,8'he4,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'h00,8'h00,8'h00,8'he4,8'he4,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'h00,8'h00,8'h00,8'h00,8'h00,8'he4,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'he4,8'h00,8'h00,8'h00,8'h00,8'h00,8'he4,8'h00,8'h00,8'h62,8'h62,8'h62}};

const logic[0:15][0:15][7:0] ai_car_yellow = {
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'hf8,8'hff,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hf8,8'hff,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hff,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hff,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hff,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hff,8'h00,8'h00,8'h00,8'hf8,8'hf8,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h91,8'h00,8'h00,8'h00,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'hf8,8'hf8,8'hf8,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'hf8,8'hf8,8'hf8,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'hf8,8'hf8,8'hf8,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'hf8,8'hf8,8'hf8,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hf8,8'h00,8'h00,8'h00,8'hf8,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62}};


const logic [0:31][0:127][7:0]  background = {
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h0c,8'h0c,8'h10,8'h34,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h30,8'h04,8'h04,8'h04,8'h04,8'h04,8'h2c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h74,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h0c,8'h04,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h78,8'h78,8'h78,8'h0c,8'h00,8'h04,8'h04,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h0c,8'h04,8'h04,8'h2c,8'h04,8'h0c,8'h04,8'h04,8'h00,8'h00,8'h78,8'h34,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h04,8'h30,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h0c,8'h00,8'h00,8'h0c,8'h00,8'h74,8'h30,8'h00,8'h00,8'h00,8'h10,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h74,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hbb,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h10,8'h0c,8'h99,8'h0c,8'h34,8'h0c,8'h78,8'h10,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h0c,8'hbe,8'h78,8'h79,8'h0c,8'h78,8'h04,8'h00,8'h00,8'h04,8'h74,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h9d,8'h9a,8'h2d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h99,8'h0c,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h7c,8'h00,8'h04,8'h30,8'h00,8'h00,8'h04,8'h30,8'h00,8'h04,8'h0c,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h10,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h04,8'h04,8'hbe,8'h00,8'h04,8'h04,8'h00,8'h00,8'h79,8'h38,8'h78,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h74,8'h78,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h30,8'h34,8'h00,8'h30,8'h04,8'h0c,8'h00,8'h30,8'h10,8'h78,8'h78,8'h78,8'h04,8'h2c,8'h04,8'h0c,8'h00,8'h78,8'h34,8'h10,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h2d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h0c,8'h04,8'h34,8'h0c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hbe,8'h9a,8'h04,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hbe,8'h04,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h04,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hbb,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h10,8'h30,8'h78,8'h78,8'h78,8'h34,8'h30,8'h78,8'h78,8'h30,8'h34,8'h78,8'h30,8'h74,8'h78,8'h78,8'h0c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h34,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h30,8'h34,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h2c,8'h2d,8'h00,8'h00,8'h2c,8'h78,8'h74,8'h2d,8'h00,8'h00,8'h04,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h74,8'h30,8'h30,8'h0c,8'h34,8'h78,8'h78,8'h70,8'h75,8'h00,8'h74,8'h38,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hbe,8'h9a,8'h24,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h9e,8'h04,8'h30,8'h78,8'h78,8'h78,8'h78,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h74,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h74,8'h74,8'h78,8'h78,8'h34,8'h38,8'h78,8'h74,8'h78,8'h78,8'h78,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h79,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h10,8'h30,8'h78,8'h78,8'h78,8'h78,8'h71,8'h2c,8'h00,8'h00,8'h74,8'h78,8'h75,8'h31,8'h04,8'h00,8'h0c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h00,8'h2c,8'h74,8'h0c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h0c,8'h31,8'h04,8'h00,8'h04,8'h78,8'h74,8'h2c,8'h04,8'h00,8'h04,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h04,8'h34,8'h30,8'h04,8'h00,8'h78,8'h74,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h79,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h78,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hbf,8'hba,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h34,8'h74,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h9d,8'h9a,8'h2d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h99,8'h0c,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h0c,8'h04,8'h04,8'h04,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h10,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h04,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h34,8'h78,8'h78,8'h78,8'h34,8'h00,8'h30,8'h34,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h38,8'h04,8'h04,8'h04,8'h9a,8'h00,8'h04,8'h00,8'h00,8'h00,8'h0c,8'h78,8'h78,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h70,8'h04,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h04,8'h04,8'h00,8'h0c,8'h04,8'h78,8'h10,8'h00,8'h00,8'h04,8'h34,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h0c,8'h0c,8'h9a,8'h0c,8'h0c,8'h0c,8'h34,8'h30,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h9e,8'h9a,8'h24,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h9e,8'h04,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h74,8'h75,8'h78,8'h0c,8'h74,8'h74,8'h0c,8'h04,8'h00,8'h04,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h74,8'h00,8'h30,8'h04,8'h04,8'h04,8'h0c,8'h04,8'h00,8'h04,8'h30,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h00,8'h2c,8'h70,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h78,8'h78,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h2c,8'h30,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h10,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h38,8'h0c,8'h30,8'h00,8'h74,8'h04,8'h2c,8'h00,8'h79,8'h0c,8'h78,8'h78,8'h78,8'h00,8'h00,8'h00,8'h00,8'h04,8'h30,8'h34,8'h04,8'h78,8'h78,8'h78},
	{8'h38,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h38,8'h38,8'h38,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hbe,8'h96,8'h04,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hbe,8'h04,8'h30,8'h38,8'h38,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h10,8'h04,8'h04,8'h04,8'h0c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h10,8'h78,8'h10,8'h78,8'h10,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78}};

const logic[0:15][0:15][7:0] finish_line = {
	{8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00, 8'hFF},
	{8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF, 8'h00},
	{8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00, 8'hFF},
	{8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF, 8'h00},
	{8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00, 8'hFF},
	{8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF, 8'h00},
	{8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00, 8'hFF},
	{8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF, 8'h00},
	{8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00, 8'hFF},
	{8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF, 8'h00},
	{8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00, 8'hFF},
	{8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF, 8'h00},
	{8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00, 8'hFF},
	{8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF, 8'h00},
	{8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00, 8'hFF},
	{8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF,8'h00,8'hFF, 8'h00}};

localparam logic[7:0] MASK_VALUE = 8'h62;
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
			RGBout <= 1'b0;
	end
	
	else begin
	//// --------------
	//// sprite priority
	//// --------------
		if(player_car_color != MASK_VALUE) begin
			RGBout <= player_car_color;
		end
		else if(ai_car_color != MASK_VALUE) begin
			RGBout <= ai_car_color;
		end
		else if(fl_color != MASK_VALUE) begin
			RGBout <= fl_color;
		end
		else if(bg_color != MASK_VALUE) begin
			RGBout <= bg_color;
		end
		else begin
			RGBout <= 8'b0000_0000;
		end
		
	//// --------------
	//// collisions
	//// --------------
		if(requested_x == 1 && requested_y == 1) begin
			collisions[0] <= 0;
			collisions[1] <= 0;
		end
		else begin
			if(player_car_color != MASK_VALUE) begin
				if(ai_car_color != MASK_VALUE) begin
					collisions[0] <= 1'd1;
				end	
				if(fl_color != MASK_VALUE) begin
					collisions[1] <= 1'd1;
				end
			end
		end
	end
end

always begin
	integer i,j;
	for (i=0; i<16; i=i+1) for (j=0; j<16; j=j+1) out_ai_car_red[j*16+i] = ai_car_red[j][i];
	for (i=0; i<16; i=i+1) for (j=0; j<16; j=j+1) out_ai_car_yellow[j*16+i] = ai_car_yellow[j][i];
	for (i=0; i<16; i=i+1) for (j=0; j<16; j=j+1) out_car1[j*16+i] = car1[j][i];
	for (i=0; i<16; i=i+1) for (j=0; j<16; j=j+1) out_car2[j*16+i] = car2[j][i];
	for (i=0; i<16; i=i+1) for (j=0; j<16; j=j+1) out_car3[j*16+i] = car3[j][i];
	for (i=0; i<128; i=i+1) for (j=0; j<32; j=j+1) out_background[j*128+i] = background[j][i];
	for (i=0; i<16; i=i+1) for (j=0; j<16; j=j+1) out_finish_line[j*16+i] = finish_line[j][i];
end

endmodule
