module	sprite_storage	(	
//		--------	Clock Input	 	
					input		logic	clk,
					input		logic	resetN,
					input    logic frame_start,
					input    int sprite_number,
					input    int requested_x,
					input    int requested_y,
					input    int x_offset,
					input    int y_offset,
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
);
localparam  int OBJECT_NUMBER_OF_Y_BITS = 7;  // 2^5 = 32 
localparam  int OBJECT_NUMBER_OF_X_BITS = 7;  // 2^6 = 64 
localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;
localparam  int OBJECT_HEIGHT_Y_DIVIDER = OBJECT_NUMBER_OF_Y_BITS - 2; //how many pixel bits are in every collision pixel
localparam  int OBJECT_WIDTH_X_DIVIDER =  OBJECT_NUMBER_OF_X_BITS - 2;
logic [0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] [7:0] object_colors = {
{8'h21, 8'h21, 8'h62, 8'h62, 8'h22, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h22, 8'h22, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h62, 8'h61, 8'h62, 8'h62, 8'h61, 8'h62, 8'h21, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h62, 8'h21, 8'h22, 8'h22, 8'h62, 8'h62, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h62, 8'h21, 8'h22, 8'h22}, 
{8'h62, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h62, 8'h21, 8'h22, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h21, 8'h62, 8'h22, 8'h62, 8'h62, 8'h21, 8'h62, 8'h61, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h21, 8'h21, 8'h61, 8'h62, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h62, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h62, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h62, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h22, 8'h22, 8'h22, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h62, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h22, 8'h21, 8'h21, 8'h22, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h21, 8'h22, 8'h61, 8'h61, 8'h21, 8'h62, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h22, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h22}, 
{8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hAD, 8'hAD, 8'h85, 8'h60, 8'h60, 8'h61, 8'h60, 8'h85, 8'hCD, 8'hA5, 8'hCD, 8'h85, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h22, 8'h22, 8'h21, 8'h21, 8'h61, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22, 8'h22, 8'h21, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h81, 8'hA5, 8'hCD, 8'hFA, 8'hFF, 8'hFF, 8'hAD, 8'hA5, 8'hA5, 8'hAD, 8'hA5, 8'hCD, 8'h60, 8'h80, 8'hA4, 8'h60, 8'h20, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h21, 8'h21, 8'h62, 8'h21, 8'h66, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h65, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h21, 8'h21, 8'h01, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h01, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h22}, 
{8'h61, 8'h61, 8'h81, 8'hA5, 8'hC5, 8'hC4, 8'hCD, 8'hAC, 8'hAD, 8'h20, 8'h60, 8'h60, 8'h20, 8'h60, 8'hFA, 8'hCD, 8'hA4, 8'hA5, 8'h60, 8'h20, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h85, 8'h21, 8'h21, 8'h85, 8'hFB, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h01, 8'h25, 8'h01, 8'h01, 8'h01, 8'h01, 8'h05, 8'h01, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h20, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h20, 8'h61, 8'h20, 8'h61, 8'h65, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'hFF, 8'h65, 8'h22}, 
{8'h61, 8'h61, 8'h81, 8'hA5, 8'hC4, 8'hC4, 8'hCC, 8'hA4, 8'h60, 8'h20, 8'hAC, 8'hFF, 8'hFF, 8'h20, 8'h60, 8'hA4, 8'hCC, 8'hA5, 8'h60, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'hFB, 8'hA5, 8'hA5, 8'h85, 8'hB1, 8'hFB, 8'hFF, 8'hFF, 8'hFB, 8'hB1, 8'hAD, 8'hAD, 8'hFB, 8'h85, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h81, 8'h81, 8'hAD, 8'hAD, 8'h8D, 8'hAD, 8'hAD, 8'h85, 8'hAD, 8'hA5, 8'hA5, 8'hAD, 8'hA5, 8'hA5, 8'hA5, 8'h85, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h26, 8'h97, 8'hBB, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'hBB, 8'h9B, 8'hBB, 8'h97, 8'hBB, 8'h9B, 8'h9B, 8'hBB, 8'hB7, 8'h21, 8'h22, 8'h22, 8'h21, 8'h21, 8'h65, 8'hD6, 8'hFA, 8'hFA, 8'hFA, 8'hFB, 8'hFA, 8'hFA, 8'hFB, 8'hFB, 8'hFB, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hD6, 8'h65, 8'h21, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'hFF, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h81, 8'hC5, 8'hE4, 8'hE4, 8'hC4, 8'h80, 8'h60, 8'h60, 8'hAC, 8'hAC, 8'hAD, 8'h20, 8'h60, 8'hAC, 8'hA4, 8'hA4, 8'h60, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'hFB, 8'hAD, 8'hA4, 8'hAD, 8'h60, 8'h20, 8'hAD, 8'hAD, 8'h84, 8'h60, 8'h60, 8'hAD, 8'hAD, 8'hFF, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h85, 8'hCD, 8'hFA, 8'hFF, 8'hFF, 8'hFF, 8'hD1, 8'h60, 8'h60, 8'h60, 8'h80, 8'hA4, 8'h60, 8'hA4, 8'hA4, 8'h80, 8'h61, 8'h21, 8'h21, 8'h21, 8'h01, 8'h97, 8'hBF, 8'hBF, 8'hBF, 8'hDF, 8'hDF, 8'h76, 8'h04, 8'h05, 8'h05, 8'h0D, 8'h9A, 8'h0D, 8'h7A, 8'h9B, 8'h01, 8'h21, 8'h21, 8'h22, 8'h21, 8'h65, 8'hD6, 8'hFF, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'hB1, 8'h20, 8'h20, 8'h20, 8'h20, 8'hFA, 8'h20, 8'hFE, 8'hFA, 8'h20, 8'h20, 8'h61, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'hFF, 8'h20, 8'h22}, 
{8'h61, 8'h61, 8'h81, 8'hA5, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'h60, 8'h80, 8'hA4, 8'hCD, 8'hA4, 8'h60, 8'h60, 8'hAC, 8'hA4, 8'hA5, 8'h60, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'hFF, 8'hA5, 8'hA5, 8'h60, 8'h20, 8'h20, 8'hAC, 8'hA4, 8'hA4, 8'h60, 8'h60, 8'hAD, 8'h8D, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'hFB, 8'hFA, 8'hCD, 8'hA4, 8'hAD, 8'h20, 8'h20, 8'hA4, 8'hA4, 8'hCC, 8'hAC, 8'h60, 8'h60, 8'hAC, 8'hA4, 8'h60, 8'h61, 8'h61, 8'h21, 8'h21, 8'h01, 8'hDF, 8'hBF, 8'h7F, 8'h7F, 8'h9A, 8'h04, 8'h00, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h04, 8'h05, 8'h9A, 8'hBB, 8'h01, 8'h01, 8'h21, 8'h21, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'hF9, 8'hF9, 8'hFA, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'h20, 8'h20, 8'hFA, 8'hFA, 8'h20, 8'h20, 8'h61, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h60, 8'h80, 8'hA0, 8'hA0, 8'hA0, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h60, 8'h60, 8'h80, 8'h20, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h65, 8'hFA, 8'hFA, 8'hFA, 8'hFB, 8'h20, 8'h21, 8'h21, 8'h21, 8'h61, 8'hFF, 8'hAD, 8'hAD, 8'h60, 8'h20, 8'h60, 8'hA4, 8'hAD, 8'hAD, 8'h20, 8'h60, 8'hAD, 8'h8D, 8'hFF, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h60, 8'hCD, 8'hCC, 8'hC4, 8'hCC, 8'hA4, 8'h20, 8'h20, 8'hA4, 8'hCC, 8'hA4, 8'hA4, 8'h60, 8'h60, 8'hAC, 8'hA4, 8'h60, 8'h61, 8'h61, 8'h21, 8'h21, 8'h05, 8'h7B, 8'h7F, 8'h3F, 8'h7F, 8'h7A, 8'h04, 8'h04, 8'hBF, 8'h7A, 8'h9F, 8'h9A, 8'h04, 8'h04, 8'h9B, 8'h9B, 8'h01, 8'h01, 8'h21, 8'h21, 8'h21, 8'h20, 8'hFA, 8'hF9, 8'hF9, 8'hFE, 8'hFA, 8'h00, 8'h00, 8'hFE, 8'hFE, 8'hF9, 8'hFA, 8'h00, 8'h20, 8'hFE, 8'hFA, 8'h20, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h86, 8'hFF, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'h80, 8'h80, 8'h80, 8'h80, 8'h60, 8'h20, 8'h20, 8'h20, 8'h20, 8'h64, 8'h60, 8'h60, 8'h60, 8'h20, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h21, 8'h61, 8'h20, 8'hFE, 8'hFA, 8'hFA, 8'hF6, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'hFF, 8'hAD, 8'hA5, 8'hAD, 8'h60, 8'h20, 8'hAD, 8'hAD, 8'h84, 8'h60, 8'h60, 8'hA4, 8'h8D, 8'hFF, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hC4, 8'hC4, 8'hE4, 8'hC4, 8'h60, 8'h60, 8'hA4, 8'hCC, 8'hA4, 8'hA4, 8'h80, 8'h60, 8'hAC, 8'hA4, 8'h60, 8'h61, 8'h61, 8'h21, 8'h21, 8'h05, 8'h7B, 8'h7F, 8'h3E, 8'h3F, 8'h7E, 8'h0D, 8'h04, 8'h76, 8'h9A, 8'h9A, 8'h7A, 8'h0D, 8'h04, 8'h9A, 8'h9A, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h65, 8'hFA, 8'hFA, 8'hF9, 8'hF9, 8'hF9, 8'h64, 8'h20, 8'hD6, 8'hFA, 8'hFA, 8'hFA, 8'h20, 8'h00, 8'hFE, 8'hFA, 8'h20, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h65, 8'h22}, 
{8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'h60, 8'h20, 8'h20, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h20, 8'h20, 8'h20, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h60, 8'hFA, 8'hFA, 8'hFA, 8'h64, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'hFF, 8'hA5, 8'hAD, 8'h8D, 8'hAD, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'hAD, 8'hAD, 8'hAD, 8'hFF, 8'h85, 8'h21, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hCD, 8'hC4, 8'hC4, 8'hC4, 8'h84, 8'h60, 8'h60, 8'h80, 8'h60, 8'h80, 8'h84, 8'h60, 8'hAC, 8'hA4, 8'h60, 8'h21, 8'h21, 8'h21, 8'h21, 8'h01, 8'h7B, 8'h9F, 8'h7F, 8'h3E, 8'h7E, 8'h36, 8'h0C, 8'h04, 8'h0C, 8'h0C, 8'h0D, 8'h35, 8'h0D, 8'h9A, 8'h9A, 8'h01, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'hD6, 8'hFE, 8'hF9, 8'hF9, 8'hFE, 8'hD5, 8'h20, 8'h20, 8'h20, 8'h00, 8'h00, 8'hDA, 8'h64, 8'hFA, 8'hFA, 8'h20, 8'h20, 8'h61, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h00, 8'h20, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h60, 8'hFA, 8'hFA, 8'hFA, 8'h20, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h85, 8'h21, 8'h21, 8'h65, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h60, 8'h84, 8'hA4, 8'hA4, 8'hA4, 8'hAD, 8'h8C, 8'hAC, 8'hAC, 8'hAC, 8'hAD, 8'hAD, 8'h84, 8'hAD, 8'hAD, 8'h85, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h05, 8'h76, 8'h9B, 8'h7A, 8'h9E, 8'h9E, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'hBE, 8'h9A, 8'h9A, 8'hBB, 8'h97, 8'h21, 8'h21, 8'h21, 8'h61, 8'h20, 8'h64, 8'hD5, 8'hFA, 8'hFA, 8'hFA, 8'hFE, 8'hDA, 8'hDA, 8'hFA, 8'hFA, 8'hFE, 8'hFE, 8'hDA, 8'hFA, 8'hFF, 8'hD6, 8'h85, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h22}, 
{8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'hFB, 8'hF6, 8'h85, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h66, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h20, 8'h20, 8'h60, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h60, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h05, 8'h04, 8'h04, 8'h04, 8'h04, 8'h00, 8'h00, 8'h00, 8'h04, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h00, 8'h20, 8'h00, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hD7, 8'h85, 8'h20, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h20, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h20, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h62, 8'h62, 8'h22, 8'h61, 8'h21, 8'h21, 8'h22}, 
{8'h21, 8'h21, 8'h62, 8'h22, 8'h21, 8'h22, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h22, 8'h62, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h62, 8'h22, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h22, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h22, 8'h22, 8'h62, 8'h61, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h21, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h65, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h22, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h01, 8'h21, 8'h01, 8'h21, 8'h21, 8'h21, 8'h22, 8'h62, 8'h21, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h62, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hA5, 8'h60, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h66, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h66, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h21, 8'h21, 8'h01, 8'h01, 8'h21, 8'h01, 8'h01, 8'h25, 8'h01, 8'h26, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h60, 8'hAD, 8'hA5, 8'hA5, 8'h60, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h25, 8'hBB, 8'h9B, 8'h9A, 8'hBB, 8'h01, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h60, 8'h85, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h01, 8'h01, 8'h05, 8'h01, 8'h01, 8'h05, 8'h01, 8'h01, 8'h01, 8'h05, 8'h01, 8'h05, 8'h01, 8'h25, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h20, 8'h61, 8'h20, 8'h61, 8'h20, 8'h65, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h22}, 
{8'h61, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'hCD, 8'hFA, 8'hCC, 8'hCD, 8'hA4, 8'h80, 8'h60, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h01, 8'h9B, 8'h7B, 8'h9F, 8'h9B, 8'h01, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h81, 8'h85, 8'hAD, 8'hAD, 8'h8D, 8'h8D, 8'h85, 8'hAD, 8'hAD, 8'hAD, 8'h85, 8'hA5, 8'hA5, 8'hAD, 8'h85, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h01, 8'h2E, 8'h97, 8'h9B, 8'h97, 8'hBB, 8'h97, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'hBB, 8'h9B, 8'hBB, 8'hBB, 8'hB7, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h20, 8'h85, 8'hF6, 8'hFA, 8'hFA, 8'hFB, 8'hFB, 8'hFA, 8'hFF, 8'hFA, 8'hFB, 8'hFB, 8'hFA, 8'hFA, 8'hFB, 8'hF7, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'hAD, 8'hFA, 8'hCD, 8'hA4, 8'hCC, 8'hC4, 8'hC4, 8'h80, 8'h60, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h22, 8'h62, 8'h21, 8'h21, 8'h06, 8'h9B, 8'h7B, 8'h7B, 8'h05, 8'h01, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h81, 8'hA5, 8'hCD, 8'hFA, 8'hFF, 8'hFF, 8'h20, 8'h20, 8'h60, 8'hFF, 8'h60, 8'hAD, 8'hA4, 8'h80, 8'hA5, 8'h60, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h01, 8'h06, 8'h77, 8'h9F, 8'hBF, 8'hFF, 8'hFF, 8'h04, 8'h00, 8'h04, 8'hFF, 8'h05, 8'h9A, 8'h9B, 8'h0D, 8'h9B, 8'h01, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h85, 8'hD6, 8'hFE, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h20, 8'h00, 8'hFF, 8'h20, 8'hFA, 8'hFE, 8'h20, 8'hF6, 8'h20, 8'h20, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h65, 8'h22}, 
{8'h22, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hAD, 8'h20, 8'h60, 8'hA4, 8'hCC, 8'hC4, 8'hC4, 8'hA4, 8'h80, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h01, 8'h01, 8'h9B, 8'h9F, 8'h9B, 8'h01, 8'h01, 8'h21, 8'h62, 8'h62, 8'h21, 8'h22, 8'h22, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h81, 8'hC5, 8'hC5, 8'hC4, 8'hA4, 8'h20, 8'h00, 8'h20, 8'hFF, 8'hFF, 8'h60, 8'h20, 8'h60, 8'hA4, 8'h80, 8'hA4, 8'h60, 8'h61, 8'h61, 8'h21, 8'h22, 8'h21, 8'h01, 8'h7B, 8'h7F, 8'h3F, 8'h3A, 8'h04, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h04, 8'h00, 8'h04, 8'h7A, 8'h0D, 8'h9B, 8'h01, 8'h01, 8'h21, 8'h21, 8'h21, 8'h61, 8'hF6, 8'hFA, 8'hF9, 8'hFA, 8'h20, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h20, 8'h00, 8'h20, 8'hFA, 8'h20, 8'hFE, 8'h00, 8'h65, 8'h61, 8'h21, 8'h61, 8'h21, 8'h22, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22}, 
{8'h22, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'hAD, 8'hFF, 8'h60, 8'h60, 8'h60, 8'hA4, 8'hC4, 8'hC4, 8'hC4, 8'hA5, 8'hA5, 8'h81, 8'h61, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h01, 8'hBB, 8'h97, 8'h05, 8'h01, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'hC5, 8'hC4, 8'hC4, 8'hCC, 8'h20, 8'h20, 8'h20, 8'h8D, 8'hAD, 8'hAD, 8'h20, 8'h60, 8'hAC, 8'hA4, 8'hAD, 8'h60, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h05, 8'h7B, 8'h3F, 8'h3F, 8'h7F, 8'h00, 8'h00, 8'h00, 8'hBA, 8'h9A, 8'h9A, 8'h00, 8'h04, 8'h9A, 8'h9A, 8'h9B, 8'h01, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'hFA, 8'hFA, 8'hF9, 8'hFA, 8'h00, 8'h00, 8'h00, 8'hFE, 8'hFA, 8'hFA, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'h20, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h22}, 
{8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'hAD, 8'hFF, 8'hAD, 8'h84, 8'h60, 8'h60, 8'h80, 8'hC4, 8'hC4, 8'hC4, 8'hA5, 8'hA5, 8'h81, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'hB7, 8'h05, 8'h01, 8'h21, 8'h22, 8'h61, 8'h61, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'hC5, 8'hC4, 8'hC4, 8'hC4, 8'h20, 8'h20, 8'h20, 8'hAC, 8'hAC, 8'hAC, 8'h60, 8'h60, 8'hA4, 8'hA4, 8'hAD, 8'h60, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h01, 8'h9F, 8'h3F, 8'h3F, 8'h7F, 8'h04, 8'h00, 8'h04, 8'h9A, 8'h9A, 8'h9A, 8'h04, 8'h00, 8'h9F, 8'h7A, 8'h9B, 8'h01, 8'h01, 8'h21, 8'h21, 8'h61, 8'h60, 8'hFA, 8'hF9, 8'hF9, 8'hFE, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFE, 8'h00, 8'h20, 8'hFA, 8'hFA, 8'hFA, 8'h20, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h22}, 
{8'h62, 8'h21, 8'h61, 8'h61, 8'hA5, 8'hAD, 8'hFF, 8'h20, 8'h60, 8'h84, 8'hAD, 8'hA4, 8'hA4, 8'h80, 8'hA0, 8'h80, 8'h80, 8'h60, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h22, 8'h01, 8'h26, 8'h01, 8'h21, 8'h22, 8'h21, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h65, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h66, 8'h21, 8'h21, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hC4, 8'hC4, 8'hA4, 8'h60, 8'h20, 8'h60, 8'hA4, 8'hAC, 8'hA4, 8'h60, 8'h60, 8'hA4, 8'h80, 8'hA5, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h05, 8'h7B, 8'h7F, 8'h3E, 8'h3E, 8'h0C, 8'h00, 8'h04, 8'h9A, 8'h9F, 8'h7A, 8'h04, 8'h0D, 8'h7A, 8'h0D, 8'h9B, 8'h01, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'hF6, 8'hFE, 8'hF9, 8'hF9, 8'h24, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'h20, 8'h20, 8'hFA, 8'h20, 8'hFE, 8'h00, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h61, 8'h61, 8'hA5, 8'hFB, 8'hAD, 8'h60, 8'h20, 8'h60, 8'h84, 8'h80, 8'h80, 8'h80, 8'h80, 8'h80, 8'h20, 8'h20, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h22, 8'h21, 8'h22, 8'h22, 8'h21, 8'h62, 8'h21, 8'h62, 8'h22, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'hFF, 8'hFF, 8'hFF, 8'hFB, 8'h65, 8'h21, 8'h21, 8'h20, 8'h65, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h65, 8'h21, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h80, 8'hA4, 8'hC4, 8'hCC, 8'hA4, 8'h60, 8'h20, 8'h60, 8'h60, 8'h60, 8'h60, 8'hA4, 8'hAC, 8'h60, 8'hAD, 8'h60, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h01, 8'h05, 8'h36, 8'h7F, 8'h7F, 8'h7A, 8'h04, 8'h04, 8'h04, 8'h04, 8'h0D, 8'h04, 8'h9A, 8'h9A, 8'h0D, 8'h7A, 8'h05, 8'h21, 8'h21, 8'h21, 8'h21, 8'h20, 8'h60, 8'hD5, 8'hFE, 8'hFE, 8'hD5, 8'h24, 8'h00, 8'h20, 8'h20, 8'h00, 8'h00, 8'hFA, 8'hFE, 8'h20, 8'hFA, 8'h20, 8'h20, 8'h21, 8'h62, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h65, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'hA5, 8'hFF, 8'hA4, 8'hCC, 8'hA4, 8'h60, 8'h60, 8'h80, 8'h60, 8'h60, 8'h60, 8'h60, 8'h20, 8'h20, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h62, 8'h22, 8'h22, 8'h21, 8'h61, 8'h61, 8'hFF, 8'hA5, 8'hAD, 8'h84, 8'hD2, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hFF, 8'hFF, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h60, 8'h60, 8'hA4, 8'hAC, 8'hAD, 8'h84, 8'hAD, 8'h8D, 8'h8C, 8'hAC, 8'h84, 8'hAD, 8'hAD, 8'h84, 8'hAD, 8'h85, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h01, 8'h01, 8'h05, 8'h7B, 8'h7A, 8'hBF, 8'h9A, 8'hBA, 8'hBA, 8'hBA, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h76, 8'hBF, 8'h96, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h20, 8'h64, 8'hFA, 8'hDA, 8'hFE, 8'hFA, 8'hFE, 8'hFA, 8'hFA, 8'hFA, 8'hFE, 8'hFA, 8'hFA, 8'hFA, 8'hFE, 8'hD6, 8'h65, 8'h21, 8'h21, 8'h22, 8'h21, 8'h62, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'hA5, 8'hA4, 8'hC4, 8'hC4, 8'hC4, 8'hA4, 8'h80, 8'h84, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'hFF, 8'hAD, 8'hC4, 8'hC4, 8'hCC, 8'h84, 8'h60, 8'h00, 8'h00, 8'hD6, 8'h20, 8'h00, 8'hFA, 8'hFA, 8'hFF, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h00, 8'h00, 8'h00, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h00, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h00, 8'h00, 8'h04, 8'h00, 8'h00, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h00, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h00, 8'h21, 8'h62, 8'h62, 8'h22, 8'h61, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'hA5, 8'hCD, 8'hC4, 8'hE4, 8'hC4, 8'hA4, 8'hA4, 8'h60, 8'h20, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h62, 8'h61, 8'h62, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'hFB, 8'hA5, 8'hC4, 8'hC4, 8'hC4, 8'h60, 8'h20, 8'hDA, 8'hFE, 8'hFE, 8'h00, 8'h00, 8'hFE, 8'hFA, 8'hFF, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h20, 8'h20, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h81, 8'hA5, 8'hC5, 8'hC4, 8'hC4, 8'hCD, 8'hA4, 8'h60, 8'h20, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'hFF, 8'hA4, 8'hC4, 8'hC4, 8'hA4, 8'h60, 8'h00, 8'hDE, 8'hDE, 8'hDE, 8'h00, 8'h00, 8'hDE, 8'hDE, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h81, 8'hA5, 8'hC5, 8'hA5, 8'h60, 8'h20, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'hFF, 8'hAD, 8'hC4, 8'hC4, 8'hC4, 8'h60, 8'h00, 8'hBA, 8'hBA, 8'hBA, 8'h00, 8'h00, 8'h9A, 8'hBA, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h01, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h61, 8'h21, 8'h21, 8'h61, 8'hFF, 8'hAD, 8'hA4, 8'hCC, 8'hC4, 8'hA4, 8'h20, 8'h00, 8'h04, 8'h96, 8'h04, 8'h04, 8'h9A, 8'h9A, 8'hFF, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h22, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h20, 8'hFF, 8'hAD, 8'hA4, 8'hA4, 8'hD1, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hBA, 8'h9A, 8'hBA, 8'hFF, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h22, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h22, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h22}, 
{8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'h20, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h65, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h20, 8'h00, 8'h00, 8'h00, 8'h04, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h25, 8'h21, 8'h22, 8'h22, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h62, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h21, 8'h62, 8'h21, 8'h22, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h20, 8'hFF, 8'hFF, 8'h22}, 
{8'h62, 8'h62, 8'h21, 8'h21, 8'h22, 8'h22, 8'h61, 8'h61, 8'h61, 8'h60, 8'hA5, 8'hA5, 8'hAD, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h01, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h01, 8'h21, 8'h21, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'hFF, 8'h21, 8'h22}, 
{8'h22, 8'h22, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h60, 8'hCD, 8'hA4, 8'hCD, 8'hA4, 8'h80, 8'h60, 8'h60, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h60, 8'h61, 8'h61, 8'h60, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h22, 8'h22, 8'h22, 8'h21, 8'h25, 8'h01, 8'h21, 8'h01, 8'h25, 8'h05, 8'h01, 8'h05, 8'h05, 8'h01, 8'h05, 8'h01, 8'h21, 8'h01, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h65, 8'h20, 8'h20, 8'h20, 8'h65, 8'h61, 8'h20, 8'h20, 8'h20, 8'h61, 8'h20, 8'h20, 8'h65, 8'h20, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'hFF, 8'h21, 8'h22}, 
{8'h22, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'hAD, 8'hA4, 8'hFA, 8'hA4, 8'hCD, 8'hA4, 8'hCD, 8'h60, 8'h60, 8'h60, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h61, 8'h62, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hAD, 8'h60, 8'h60, 8'h60, 8'hA5, 8'h85, 8'hAD, 8'hAD, 8'hA5, 8'hA5, 8'hAD, 8'h60, 8'h60, 8'h80, 8'h85, 8'h61, 8'h61, 8'h61, 8'h22, 8'h22, 8'h21, 8'h26, 8'h72, 8'h05, 8'h01, 8'h05, 8'h77, 8'h9B, 8'hBB, 8'h9B, 8'h9B, 8'hBB, 8'h97, 8'h01, 8'h00, 8'h05, 8'hB7, 8'h21, 8'h21, 8'h22, 8'h21, 8'h21, 8'h65, 8'hD6, 8'h20, 8'h20, 8'h20, 8'hFA, 8'hFA, 8'hFB, 8'hFF, 8'hFA, 8'hFA, 8'hFA, 8'h20, 8'h20, 8'h20, 8'hD7, 8'h61, 8'h21, 8'h62, 8'h22, 8'h62, 8'h62, 8'h21, 8'h21, 8'hFF, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h81, 8'hA5, 8'hFB, 8'h60, 8'hAC, 8'hA4, 8'hCC, 8'hC4, 8'hC4, 8'hC4, 8'hA5, 8'hA5, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hCD, 8'hFA, 8'hCD, 8'hC4, 8'hA4, 8'hCC, 8'hAD, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFA, 8'hCD, 8'hA4, 8'hA4, 8'hA5, 8'h61, 8'h61, 8'h61, 8'h22, 8'h21, 8'h01, 8'h9B, 8'hBF, 8'h7F, 8'h3B, 8'h7F, 8'h7F, 8'h9F, 8'hDF, 8'hDF, 8'hDF, 8'hBF, 8'hBF, 8'h9F, 8'h7A, 8'h9B, 8'h9B, 8'h01, 8'h21, 8'h21, 8'h61, 8'h61, 8'hF6, 8'hFF, 8'hF9, 8'hFE, 8'hF9, 8'hFE, 8'hFE, 8'hFF, 8'hFE, 8'hFF, 8'hFE, 8'hFE, 8'hFE, 8'hFA, 8'hFA, 8'hFB, 8'h20, 8'h21, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h65, 8'hFB, 8'h65, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hAD, 8'hA4, 8'h60, 8'h60, 8'h60, 8'hA4, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hA5, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h62, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h62, 8'h21, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hCD, 8'hC4, 8'hE4, 8'hC4, 8'hC4, 8'hFF, 8'hFF, 8'h60, 8'hAC, 8'hAC, 8'hCD, 8'hA4, 8'h80, 8'hC4, 8'hC5, 8'h61, 8'h61, 8'h61, 8'h22, 8'h21, 8'h01, 8'h9B, 8'h7F, 8'h3F, 8'h3F, 8'h3F, 8'h7F, 8'hDF, 8'hFF, 8'h04, 8'h7A, 8'h7E, 8'h7E, 8'h7A, 8'h0D, 8'h7B, 8'h9F, 8'h01, 8'h21, 8'h21, 8'h21, 8'h60, 8'hFA, 8'hF9, 8'hF9, 8'hF9, 8'hFD, 8'hF9, 8'hFE, 8'hFF, 8'h20, 8'hF9, 8'hFE, 8'hF9, 8'hF9, 8'h20, 8'hFA, 8'hFA, 8'h60, 8'h61, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h21, 8'h65, 8'h21, 8'h22}, 
{8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h61, 8'hA5, 8'hFA, 8'hCD, 8'hA4, 8'h60, 8'h60, 8'h60, 8'h80, 8'hC4, 8'hC4, 8'hA4, 8'h60, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h21, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h22, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hC4, 8'hC4, 8'hE4, 8'hC4, 8'hC4, 8'hFE, 8'h20, 8'h20, 8'hAC, 8'hAC, 8'hC4, 8'hC4, 8'h80, 8'hC4, 8'hC5, 8'h81, 8'h61, 8'h61, 8'h21, 8'h21, 8'h01, 8'h7B, 8'h3F, 8'h1F, 8'h3F, 8'h3F, 8'h7F, 8'hDF, 8'h04, 8'h04, 8'h9A, 8'h7E, 8'h7F, 8'h7E, 8'h0D, 8'h7F, 8'h7B, 8'h01, 8'h21, 8'h21, 8'h61, 8'h20, 8'hFA, 8'hF9, 8'hF9, 8'hF9, 8'hF9, 8'hFE, 8'hFE, 8'h20, 8'h00, 8'hFE, 8'hF9, 8'hF9, 8'hF9, 8'h20, 8'hFA, 8'hFA, 8'h60, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'h21, 8'h22}, 
{8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h60, 8'hCD, 8'h84, 8'hAD, 8'hA4, 8'h60, 8'h60, 8'h80, 8'hA4, 8'hA4, 8'h80, 8'h60, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hED, 8'hC4, 8'hE4, 8'hC4, 8'hC4, 8'h60, 8'h20, 8'h60, 8'hAC, 8'hA4, 8'hA4, 8'hA4, 8'h80, 8'hC4, 8'hC5, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h01, 8'h9F, 8'h7F, 8'h3F, 8'h3E, 8'h3F, 8'h3A, 8'h0D, 8'h00, 8'h04, 8'h9A, 8'h7E, 8'h7A, 8'h7A, 8'h0D, 8'h7B, 8'h9B, 8'h05, 8'h21, 8'h21, 8'h21, 8'h60, 8'hFA, 8'hFA, 8'hF9, 8'hF9, 8'hFD, 8'hD5, 8'h64, 8'h00, 8'h20, 8'hFA, 8'hFA, 8'hFA, 8'hF9, 8'h20, 8'hF6, 8'hFF, 8'h20, 8'h21, 8'h61, 8'h61, 8'h62, 8'h21, 8'h21, 8'h61, 8'hFB, 8'h65, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'hAD, 8'h84, 8'h80, 8'hAC, 8'hA4, 8'hAD, 8'hA4, 8'hA4, 8'hAC, 8'h80, 8'h20, 8'h20, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hAD, 8'hFA, 8'hCD, 8'hC4, 8'hA4, 8'hA4, 8'hAC, 8'h60, 8'h60, 8'h60, 8'h60, 8'h80, 8'hA4, 8'hA4, 8'hA4, 8'hAD, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h01, 8'h9B, 8'hBF, 8'h7F, 8'h7E, 8'h3A, 8'h9F, 8'h76, 8'h0C, 8'h04, 8'h04, 8'h04, 8'h0D, 8'h9A, 8'h9A, 8'h9B, 8'h9B, 8'h01, 8'h01, 8'h61, 8'h21, 8'h61, 8'hF6, 8'hFF, 8'hF9, 8'hFA, 8'hF9, 8'hFE, 8'hD5, 8'h20, 8'h00, 8'h00, 8'h00, 8'h20, 8'hFA, 8'hFA, 8'hFA, 8'hFB, 8'h20, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h21, 8'h21, 8'h66, 8'h21, 8'h22}, 
{8'h62, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'hCE, 8'hFB, 8'h60, 8'h60, 8'h60, 8'h60, 8'hA4, 8'hA4, 8'h60, 8'h60, 8'h20, 8'h20, 8'h21, 8'h21, 8'h21, 8'h62, 8'h22, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h62, 8'h61, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'hAD, 8'h60, 8'h20, 8'h60, 8'hAC, 8'hAC, 8'h8C, 8'hAD, 8'h8D, 8'hAD, 8'h84, 8'h60, 8'h20, 8'h60, 8'h85, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h01, 8'h97, 8'h05, 8'h04, 8'h0D, 8'h7A, 8'hBF, 8'h9A, 8'h9A, 8'h9A, 8'hBF, 8'h76, 8'h04, 8'h00, 8'h0D, 8'h97, 8'h01, 8'h21, 8'h21, 8'h21, 8'h20, 8'h65, 8'hD6, 8'h20, 8'h00, 8'h20, 8'hDA, 8'hFE, 8'hFA, 8'hFA, 8'hFA, 8'hFA, 8'hDA, 8'h20, 8'h00, 8'h20, 8'hD6, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'hFB, 8'hAD, 8'hA4, 8'h80, 8'h60, 8'h80, 8'hA4, 8'h60, 8'h20, 8'h20, 8'h20, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h22, 8'h22, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h20, 8'h20, 8'h20, 8'h00, 8'h20, 8'h20, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h21, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h62, 8'h21, 8'h61, 8'h22}, 
{8'h22, 8'h22, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hFB, 8'hA4, 8'hCC, 8'hA4, 8'hA4, 8'hA4, 8'h84, 8'h20, 8'h20, 8'h00, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h86, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h65, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h22, 8'h61, 8'h21, 8'h21, 8'h22}, 
{8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hCD, 8'hC4, 8'hC4, 8'hC4, 8'hCD, 8'hA5, 8'h60, 8'h20, 8'h00, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h85, 8'h61, 8'h21, 8'h65, 8'h85, 8'h61, 8'h61, 8'h81, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h66, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'h80, 8'h20, 8'h20, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h22, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h22, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h85, 8'h61, 8'hFF, 8'hAD, 8'h60, 8'hAE, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22}, 
{8'h62, 8'h61, 8'h62, 8'h61, 8'h61, 8'h81, 8'hA5, 8'hC5, 8'hC5, 8'hC5, 8'hA5, 8'h60, 8'h20, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'hFF, 8'h8D, 8'h00, 8'hFF, 8'h8D, 8'h20, 8'hAE, 8'h61, 8'h86, 8'h61, 8'h61, 8'h61, 8'h61, 8'h22, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h65, 8'h20, 8'h22}, 
{8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h61, 8'h81, 8'h80, 8'h80, 8'h80, 8'h60, 8'h60, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h20, 8'h20, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'hAD, 8'hFF, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h22, 8'h22, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h22, 8'h62, 8'h61, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h22}, 
{8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h8E, 8'h61, 8'h85, 8'hFF, 8'h00, 8'hFF, 8'hFF, 8'h20, 8'hA5, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h22, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h22, 8'h22, 8'h22, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h61, 8'h21, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h62, 8'h21, 8'h22, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h22}, 
{8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h8D, 8'hFF, 8'hFF, 8'h8D, 8'hFF, 8'hFF, 8'hAD, 8'h85, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h22, 8'h22, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h25, 8'h22}, 
{8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'hA5, 8'hA5, 8'h80, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'hA5, 8'hA5, 8'h60, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'hFB, 8'hAE, 8'h60, 8'h20, 8'h20, 8'h8D, 8'hFF, 8'h20, 8'hAD, 8'h60, 8'hAD, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h62, 8'h61, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h01, 8'h25, 8'h01, 8'h21, 8'h21, 8'h01, 8'h25, 8'h25, 8'h01, 8'h26, 8'h05, 8'h01, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h65, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h20, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'hC5, 8'hC5, 8'hA4, 8'hCC, 8'hCD, 8'hA4, 8'hC4, 8'hC4, 8'hC4, 8'hC5, 8'h60, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h85, 8'h20, 8'h20, 8'hAD, 8'h85, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h20, 8'hB2, 8'hFB, 8'hFF, 8'h00, 8'h20, 8'h60, 8'hA5, 8'hA5, 8'h60, 8'hA5, 8'hA5, 8'h81, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h22, 8'h21, 8'h21, 8'h21, 8'h01, 8'hBB, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h01, 8'h97, 8'h96, 8'h05, 8'h97, 8'h97, 8'h25, 8'h01, 8'h21, 8'h21, 8'h62, 8'h62, 8'h61, 8'h21, 8'h65, 8'h00, 8'hFB, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'h20, 8'hFB, 8'hF6, 8'h65, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h22, 8'h61, 8'h61, 8'h61, 8'hC5, 8'hC4, 8'hC4, 8'hA4, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hA4, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h20, 8'hFF, 8'h85, 8'h60, 8'hAD, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h85, 8'h80, 8'h80, 8'h60, 8'hFF, 8'h20, 8'h20, 8'h60, 8'hCC, 8'hA5, 8'h60, 8'hA4, 8'hAD, 8'h85, 8'h60, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h05, 8'h97, 8'h05, 8'h96, 8'h04, 8'hFF, 8'h00, 8'h04, 8'h05, 8'h9B, 8'h9B, 8'h05, 8'h76, 8'hBF, 8'h96, 8'h01, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'hD6, 8'h20, 8'hFA, 8'h20, 8'hFF, 8'h20, 8'h00, 8'h20, 8'hFA, 8'hFA, 8'h20, 8'hFA, 8'hFE, 8'hD5, 8'h20, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h65, 8'h22}, 
{8'h61, 8'h62, 8'h22, 8'h61, 8'h61, 8'h61, 8'hC5, 8'hC4, 8'hFA, 8'hCC, 8'hA4, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h60, 8'hAD, 8'hA4, 8'hCD, 8'h20, 8'h20, 8'hFF, 8'hAD, 8'hA4, 8'hCC, 8'hA4, 8'h60, 8'h80, 8'hA4, 8'hAD, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h01, 8'h9B, 8'h7B, 8'h9F, 8'h00, 8'h00, 8'hFF, 8'h9A, 8'h7F, 8'h7E, 8'h9A, 8'h04, 8'h0D, 8'h7A, 8'h9B, 8'h01, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h20, 8'hFE, 8'hFA, 8'hFE, 8'h00, 8'h20, 8'hFF, 8'hFE, 8'hF9, 8'hF9, 8'hF9, 8'h20, 8'h20, 8'hFA, 8'hFE, 8'h20, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h65, 8'hFF, 8'h22}, 
{8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h61, 8'hA5, 8'hA5, 8'hFF, 8'h60, 8'h20, 8'h60, 8'h60, 8'h80, 8'hC4, 8'hA5, 8'h20, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'hA6, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h22, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h60, 8'hA5, 8'hA4, 8'hAC, 8'h20, 8'h20, 8'hAC, 8'hA4, 8'hC4, 8'hC4, 8'hA4, 8'h60, 8'h60, 8'hAD, 8'hAD, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h01, 8'h9B, 8'h7F, 8'h7E, 8'h04, 8'h04, 8'h9A, 8'h7A, 8'h7F, 8'h7F, 8'h7A, 8'h04, 8'h04, 8'h9A, 8'h9A, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h20, 8'hFA, 8'hFE, 8'hFA, 8'h20, 8'h00, 8'hFA, 8'hFA, 8'hF9, 8'hF9, 8'hF9, 8'h20, 8'h00, 8'hFA, 8'hFA, 8'h20, 8'h21, 8'h21, 8'h61, 8'h21, 8'h22, 8'h21, 8'h62, 8'h21, 8'h65, 8'hFF, 8'h22}, 
{8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h80, 8'hA5, 8'hAD, 8'hFF, 8'h20, 8'h20, 8'h60, 8'hA4, 8'hAC, 8'h60, 8'h60, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h60, 8'hAD, 8'hCC, 8'hAC, 8'h20, 8'h20, 8'hAD, 8'hAC, 8'hA4, 8'hC4, 8'hA4, 8'h60, 8'h60, 8'hAC, 8'hAD, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h01, 8'h9A, 8'h9F, 8'h7A, 8'h04, 8'h04, 8'h9A, 8'h9F, 8'h3E, 8'h7E, 8'h9E, 8'h04, 8'h04, 8'h9A, 8'hBB, 8'h00, 8'h01, 8'h21, 8'h21, 8'h61, 8'h20, 8'h00, 8'hFE, 8'hF9, 8'hFE, 8'h00, 8'h64, 8'hDA, 8'hFA, 8'hFA, 8'hFD, 8'hF9, 8'h20, 8'h00, 8'hFA, 8'hFA, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h22, 8'h21, 8'h62, 8'h21, 8'h65, 8'h22}, 
{8'h61, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h80, 8'hA5, 8'hAC, 8'hFE, 8'hAD, 8'hA4, 8'hCC, 8'hA4, 8'hA4, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22, 8'h21, 8'h21, 8'h61, 8'h60, 8'h84, 8'h80, 8'h84, 8'h60, 8'h84, 8'h20, 8'h60, 8'h60, 8'hAC, 8'hAD, 8'h20, 8'h60, 8'hAC, 8'h84, 8'h20, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h9A, 8'h0C, 8'h9E, 8'h04, 8'h9A, 8'h04, 8'h00, 8'h0D, 8'h9A, 8'h9E, 8'h04, 8'h0D, 8'h9A, 8'h96, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h20, 8'hD6, 8'h24, 8'hDA, 8'h64, 8'hB1, 8'h24, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'h00, 8'h20, 8'hFE, 8'hFA, 8'h20, 8'h21, 8'h21, 8'h61, 8'h62, 8'h22, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h22}, 
{8'h62, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h60, 8'hA5, 8'hAC, 8'hFE, 8'hAC, 8'hCD, 8'hA4, 8'hCC, 8'hAC, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h86, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA6, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h20, 8'h60, 8'h84, 8'hB1, 8'h64, 8'h20, 8'h20, 8'h00, 8'h20, 8'h8C, 8'h8C, 8'h60, 8'h84, 8'h8D, 8'h20, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h04, 8'h96, 8'hBA, 8'hBA, 8'h00, 8'h00, 8'h00, 8'h04, 8'hBA, 8'h9A, 8'h04, 8'h96, 8'h9A, 8'h05, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h00, 8'h24, 8'hD6, 8'hFE, 8'hB5, 8'h24, 8'h00, 8'h00, 8'h20, 8'hFA, 8'hFA, 8'h00, 8'hDA, 8'hDA, 8'h20, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h62, 8'h61, 8'h21, 8'h21, 8'h22}, 
{8'h22, 8'h62, 8'h22, 8'h61, 8'h61, 8'h61, 8'h80, 8'hA4, 8'hAC, 8'h60, 8'h20, 8'h60, 8'h80, 8'h60, 8'hA4, 8'h60, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h81, 8'hA6, 8'h61, 8'h60, 8'h60, 8'h81, 8'h85, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hFB, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h00, 8'h00, 8'h20, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h04, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h00, 8'h00, 8'h20, 8'h00, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h61, 8'hA5, 8'hC4, 8'hA4, 8'hFE, 8'h60, 8'h60, 8'h80, 8'hC4, 8'hAD, 8'hA5, 8'h20, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hAD, 8'h60, 8'h80, 8'hA5, 8'hA5, 8'h60, 8'h61, 8'h61, 8'h61, 8'hAE, 8'hA6, 8'h61, 8'h21, 8'h62, 8'h61, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'hA5, 8'hC4, 8'hC4, 8'hCC, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hA4, 8'hAD, 8'h20, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h61, 8'h21, 8'h81, 8'h60, 8'hA5, 8'hA5, 8'hA5, 8'hA5, 8'hFB, 8'h81, 8'h60, 8'h61, 8'hA5, 8'hFF, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h22}, 
{8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'hA5, 8'hC4, 8'hC4, 8'hE4, 8'hC4, 8'hE4, 8'hC4, 8'hCD, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'hFB, 8'h60, 8'hA5, 8'hFB, 8'hAD, 8'hA5, 8'h80, 8'h60, 8'hAD, 8'hA5, 8'hFF, 8'h85, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h22, 8'h62, 8'h21, 8'h61, 8'h21, 8'h22}, 
{8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'h60, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hA4, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'hAD, 8'hA4, 8'hFF, 8'hAD, 8'hFF, 8'hAD, 8'hA5, 8'hA5, 8'hA5, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h22, 8'h21, 8'h62, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h21, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h22}, 
{8'h62, 8'h21, 8'h62, 8'h61, 8'h21, 8'h61, 8'h61, 8'h60, 8'h80, 8'hA4, 8'hC4, 8'hC4, 8'hA4, 8'h80, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hCD, 8'h84, 8'hFF, 8'h20, 8'hFF, 8'h60, 8'hAD, 8'hA4, 8'hFB, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h22, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h22, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h62, 8'h21, 8'h22, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h65, 8'h22}, 
{8'h21, 8'h62, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h20, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h85, 8'hAD, 8'hFB, 8'hCD, 8'hA4, 8'hFF, 8'hAD, 8'hFF, 8'hA4, 8'hCD, 8'hA5, 8'h60, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h21, 8'h62, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h85, 8'h20, 8'h60, 8'h60, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h81, 8'h61, 8'h60, 8'hA5, 8'hFF, 8'hAC, 8'hFF, 8'hA4, 8'h80, 8'hA5, 8'hFB, 8'hCD, 8'hA5, 8'hAE, 8'h85, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h65, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h81, 8'h81, 8'hCD, 8'hFB, 8'hCD, 8'hA5, 8'h80, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h22, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'hCE, 8'h60, 8'h60, 8'hAD, 8'hA4, 8'hFF, 8'hFB, 8'h80, 8'hC5, 8'hA5, 8'h60, 8'hFB, 8'h85, 8'h21, 8'h62, 8'h61, 8'h21, 8'h62, 8'h61, 8'h62, 8'h21, 8'h21, 8'h22, 8'h61, 8'h21, 8'h65, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h22, 8'h21, 8'h21, 8'h22, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'hA5, 8'hC5, 8'hC0, 8'hED, 8'hFA, 8'hA5, 8'hA5, 8'h80, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h22, 8'h22, 8'h61, 8'h21, 8'h61, 8'h61, 8'h81, 8'hFB, 8'h85, 8'h60, 8'hA5, 8'hA5, 8'hAD, 8'hA4, 8'hCD, 8'hA4, 8'hFB, 8'hA5, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h21, 8'h61, 8'h62, 8'h22, 8'h62, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h20, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h62, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h22, 8'h21, 8'h21, 8'h65, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h62, 8'h22, 8'h62, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h81, 8'hC5, 8'hE4, 8'hC4, 8'hA4, 8'hCD, 8'hA4, 8'hCD, 8'hA5, 8'h80, 8'h60, 8'h60, 8'h81, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h81, 8'h81, 8'hAD, 8'hFF, 8'hAD, 8'hFF, 8'hAD, 8'h60, 8'h81, 8'hA5, 8'hA5, 8'hA5, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h01, 8'h26, 8'h01, 8'h01, 8'h05, 8'h01, 8'h05, 8'h25, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h66, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h62, 8'h22, 8'h62, 8'h21, 8'h21, 8'h61, 8'h22}, 
{8'h61, 8'h61, 8'h81, 8'hC5, 8'hC4, 8'hE4, 8'hCC, 8'hA4, 8'h80, 8'h60, 8'hA4, 8'hA5, 8'hA5, 8'hA5, 8'hA5, 8'h80, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'hAD, 8'h60, 8'h60, 8'h60, 8'h60, 8'hA5, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h20, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h01, 8'h05, 8'h97, 8'h9B, 8'h9B, 8'h9B, 8'hBB, 8'h9B, 8'h05, 8'h92, 8'h92, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h92, 8'hB2, 8'h21, 8'h21, 8'h62, 8'h61, 8'h62, 8'h22, 8'h22, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h22}, 
{8'h61, 8'h61, 8'h81, 8'hC5, 8'hC4, 8'hE4, 8'hA4, 8'h60, 8'h60, 8'hFE, 8'hAD, 8'hFA, 8'hAD, 8'hA5, 8'hC5, 8'hC5, 8'h80, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h22, 8'h21, 8'h62, 8'h21, 8'h8E, 8'hFF, 8'hFF, 8'h61, 8'h61, 8'h61, 8'hFF, 8'hAE, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hFB, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h21, 8'h21, 8'h01, 8'h9B, 8'hBF, 8'h9F, 8'h9F, 8'h05, 8'h05, 8'hDF, 8'hDF, 8'h04, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h65, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h22}, 
{8'h61, 8'h61, 8'h81, 8'hA5, 8'hC5, 8'hA0, 8'h60, 8'h60, 8'h60, 8'hAD, 8'hA4, 8'hA4, 8'hFE, 8'h80, 8'hC4, 8'hC4, 8'hC5, 8'hA5, 8'h81, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h86, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h86, 8'h62, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h01, 8'h7B, 8'h7F, 8'h3A, 8'h3B, 8'h0D, 8'h9A, 8'h7A, 8'h9F, 8'h76, 8'hB6, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'hB6, 8'h01, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h81, 8'hA5, 8'hCD, 8'hA4, 8'h60, 8'hAC, 8'hA4, 8'hAC, 8'h60, 8'h60, 8'h60, 8'hC4, 8'hC4, 8'hC5, 8'hA5, 8'h85, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h01, 8'h7B, 8'h3F, 8'h3F, 8'h3F, 8'h0C, 8'h9A, 8'h7F, 8'h3A, 8'h04, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h65, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h22}, 
{8'h62, 8'h61, 8'h61, 8'h61, 8'h60, 8'h80, 8'hA5, 8'hAC, 8'hA4, 8'hCC, 8'h60, 8'h60, 8'h60, 8'hCD, 8'hC4, 8'hC4, 8'hA4, 8'h80, 8'h60, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h62, 8'h61, 8'h22, 8'h22, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h05, 8'h7F, 8'h3F, 8'h3F, 8'h3F, 8'h0C, 8'h9E, 8'h3E, 8'h7F, 8'h04, 8'h96, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'hB2, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h62, 8'h22}, 
{8'h22, 8'h62, 8'h21, 8'h61, 8'h61, 8'h60, 8'h20, 8'h60, 8'h80, 8'hA4, 8'h80, 8'h80, 8'hA4, 8'hA4, 8'hC4, 8'hA4, 8'h60, 8'h20, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h05, 8'h9F, 8'h3F, 8'h3E, 8'h3E, 8'h0D, 8'h7A, 8'h7E, 8'h7F, 8'h9A, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h65, 8'h61, 8'h21, 8'h22, 8'h62, 8'h62, 8'h62, 8'h22, 8'h62, 8'h22, 8'h22, 8'h21, 8'h61, 8'h22}, 
{8'h22, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h20, 8'h20, 8'h80, 8'h80, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hA4, 8'h60, 8'h60, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'hAE, 8'h61, 8'h61, 8'h85, 8'h61, 8'h21, 8'h61, 8'h86, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h05, 8'h77, 8'h7B, 8'h7F, 8'h7E, 8'h0C, 8'h0C, 8'h7F, 8'h7A, 8'h04, 8'h95, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h91, 8'h92, 8'hB2, 8'h01, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22, 8'h62, 8'h22, 8'h62, 8'h61, 8'h21, 8'h22}, 
{8'h22, 8'h22, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h20, 8'h20, 8'h80, 8'h80, 8'hC4, 8'hC4, 8'hC4, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'hFB, 8'hAE, 8'hFF, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h01, 8'h01, 8'h05, 8'h76, 8'h9E, 8'h9A, 8'h9A, 8'h9A, 8'h9A, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h65, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h21, 8'h62, 8'h22, 8'h61, 8'h61, 8'h21, 8'h65, 8'h22}, 
{8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h20, 8'h20, 8'h80, 8'hAC, 8'hC4, 8'h60, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h21, 8'h61, 8'h61, 8'h62, 8'h22, 8'h62, 8'h61, 8'h21, 8'h61, 8'h86, 8'h21, 8'hAE, 8'h60, 8'h60, 8'hAD, 8'h8D, 8'hFF, 8'h61, 8'hFF, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h62, 8'h21, 8'h62, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h04, 8'h00, 8'h00, 8'h00, 8'h04, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h62, 8'h21, 8'h61, 8'h21, 8'h65, 8'hFF, 8'h22}, 
{8'h22, 8'h21, 8'h22, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h20, 8'h20, 8'h60, 8'hA5, 8'hA5, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'hFF, 8'h61, 8'h20, 8'hFF, 8'h8D, 8'hAD, 8'hFF, 8'h60, 8'hAD, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h86, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h22}, 
{8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h20, 8'h20, 8'h60, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'hFF, 8'hFF, 8'h20, 8'h60, 8'hFF, 8'h20, 8'hAD, 8'hFB, 8'h61, 8'h61, 8'h61, 8'h86, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h01, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'hFF, 8'h65, 8'h22}, 
{8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'hFF, 8'h61, 8'hFF, 8'h8D, 8'h60, 8'hAD, 8'hFF, 8'hAE, 8'h20, 8'hAE, 8'hFB, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h22, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h61, 8'h61, 8'h22, 8'h22, 8'h21, 8'h61, 8'h62, 8'h61, 8'h21, 8'hFF, 8'h20, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h21, 8'h21, 8'hFF, 8'h21, 8'hFF, 8'h85, 8'h60, 8'hFF, 8'h85, 8'hFF, 8'hFF, 8'h85, 8'h85, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'hFF, 8'h65, 8'h22}, 
{8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h81, 8'h81, 8'hA5, 8'hC5, 8'hC5, 8'hAD, 8'h60, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h22, 8'h22, 8'h22, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'hFF, 8'h61, 8'h60, 8'hFF, 8'h85, 8'hFF, 8'h60, 8'h85, 8'hAE, 8'hFB, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h22, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h01, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'hFF, 8'hFF, 8'h22}, 
{8'h62, 8'h62, 8'h61, 8'h61, 8'h81, 8'hA1, 8'hC5, 8'hC5, 8'hC4, 8'hCD, 8'hFA, 8'hCE, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h22, 8'h22, 8'h22, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h62, 8'h61, 8'h21, 8'h61, 8'h61, 8'hFF, 8'h8D, 8'h8D, 8'h61, 8'h85, 8'h61, 8'h60, 8'hFB, 8'hCE, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h86, 8'hFB, 8'h22}, 
{8'h62, 8'h62, 8'h61, 8'h61, 8'h81, 8'hC5, 8'hC4, 8'hC4, 8'hC4, 8'hA4, 8'hD1, 8'hFA, 8'h85, 8'h61, 8'h61, 8'h21, 8'h61, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h85, 8'h65, 8'hFB, 8'h61, 8'hFF, 8'h61, 8'hFF, 8'h61, 8'h61, 8'h61, 8'h61, 8'h86, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h22, 8'h22, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h65, 8'h22}, 
{8'h62, 8'h21, 8'h61, 8'h61, 8'hA5, 8'hC5, 8'hC4, 8'hC4, 8'hC4, 8'hCD, 8'h60, 8'hAD, 8'hA5, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h61, 8'h61, 8'h21, 8'h21, 8'hAE, 8'h21, 8'hFF, 8'h61, 8'h61, 8'h61, 8'h86, 8'h61, 8'hFF, 8'h61, 8'h61, 8'h61, 8'h61, 8'h86, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h21, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hC5, 8'hC4, 8'hC4, 8'h60, 8'h60, 8'h60, 8'hAD, 8'hAD, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h21, 8'h62, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'hFB, 8'h61, 8'h21, 8'h61, 8'h86, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h21, 8'h62, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h22, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h81, 8'hC5, 8'hA4, 8'h60, 8'h60, 8'h20, 8'h60, 8'hFA, 8'hA5, 8'hC5, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h86, 8'h21, 8'h61, 8'h61, 8'h61, 8'hFB, 8'h86, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h22, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hA5, 8'h80, 8'h60, 8'hA4, 8'hA4, 8'hAD, 8'hA4, 8'hA5, 8'hA5, 8'hAD, 8'h81, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h62, 8'h21, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h62, 8'h61, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h65, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h80, 8'h84, 8'hAC, 8'hAC, 8'hAC, 8'h60, 8'h60, 8'h60, 8'hFB, 8'hAD, 8'hA5, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h01, 8'h01, 8'h00, 8'h00, 8'h01, 8'h01, 8'h01, 8'h21, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h20, 8'h60, 8'h80, 8'h80, 8'h60, 8'h60, 8'h60, 8'hAC, 8'hFE, 8'hA5, 8'hA5, 8'h81, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h20, 8'h8D, 8'hFF, 8'h85, 8'hAD, 8'h85, 8'h20, 8'h21, 8'h21, 8'h61, 8'h21, 8'h00, 8'hFF, 8'hFF, 8'hFA, 8'hFE, 8'hFA, 8'h20, 8'h21, 8'h61, 8'h61, 8'h21, 8'h01, 8'hBB, 8'hFF, 8'h9B, 8'h9B, 8'h96, 8'h00, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h61, 8'h62, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h22}, 
{8'h22, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h20, 8'h20, 8'h80, 8'hC4, 8'h80, 8'hA4, 8'hA4, 8'hA4, 8'hAC, 8'hFF, 8'hA5, 8'hA5, 8'h60, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h20, 8'h8D, 8'hFF, 8'hAC, 8'hAD, 8'h84, 8'h20, 8'h21, 8'h21, 8'h61, 8'h61, 8'h00, 8'hFA, 8'hFF, 8'hFA, 8'hFA, 8'hFA, 8'h20, 8'h20, 8'h61, 8'h21, 8'h21, 8'h00, 8'h9A, 8'hDF, 8'h9F, 8'h9A, 8'h9A, 8'h01, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h65, 8'h22}, 
{8'h22, 8'h21, 8'h62, 8'h61, 8'h61, 8'h21, 8'h20, 8'h20, 8'h80, 8'hA0, 8'hC4, 8'hC4, 8'hC4, 8'hCC, 8'hA4, 8'hCC, 8'hC4, 8'hA5, 8'h60, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h22, 8'h62, 8'h61, 8'h62, 8'h61, 8'h21, 8'h62, 8'h62, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h20, 8'h20, 8'h60, 8'h60, 8'h60, 8'h60, 8'h20, 8'h61, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h20, 8'h20, 8'h00, 8'h20, 8'h00, 8'h61, 8'h21, 8'h21, 8'h65, 8'h00, 8'h04, 8'h04, 8'h04, 8'h0D, 8'h04, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h20, 8'h20, 8'h80, 8'h80, 8'hA0, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'h60, 8'hA5, 8'hA5, 8'h20, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h61, 8'h62, 8'h61, 8'h21, 8'h20, 8'h8D, 8'hAD, 8'hA4, 8'hAD, 8'h85, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'hFA, 8'hFA, 8'hFA, 8'hFE, 8'hDA, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'hBA, 8'hBA, 8'h9A, 8'h9A, 8'h9A, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h62, 8'h22, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h20, 8'h80, 8'h80, 8'hA0, 8'hA4, 8'hA4, 8'h60, 8'h60, 8'h60, 8'h20, 8'h20, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h22, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h20, 8'h8D, 8'hFF, 8'hAC, 8'hAD, 8'h85, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'hFB, 8'hFF, 8'hFA, 8'hFA, 8'hFA, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'hBA, 8'hDF, 8'h9A, 8'h9A, 8'hBA, 8'h00, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h20, 8'h60, 8'h60, 8'h80, 8'h60, 8'h60, 8'h60, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h20, 8'h20, 8'h20, 8'h20, 8'h60, 8'h60, 8'h20, 8'h61, 8'h61, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h00, 8'h61, 8'h21, 8'h21, 8'h25, 8'h00, 8'h00, 8'h04, 8'h04, 8'h04, 8'h04, 8'h00, 8'h25, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h20, 8'h20, 8'h60, 8'h20, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h21, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h20, 8'h8D, 8'hFF, 8'hAC, 8'hAD, 8'h85, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h20, 8'hFA, 8'hFF, 8'hFE, 8'hFA, 8'hFA, 8'h20, 8'h21, 8'h21, 8'h21, 8'h01, 8'h00, 8'hBA, 8'hDF, 8'h9A, 8'h9A, 8'hBA, 8'h01, 8'h01, 8'h21, 8'h61, 8'h61, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h22, 8'h62, 8'h61, 8'h22}, 
{8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h20, 8'h20, 8'h20, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h21, 8'h61, 8'h21, 8'h20, 8'h8D, 8'hFF, 8'h8D, 8'hAD, 8'h85, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'hFA, 8'hFF, 8'hFA, 8'hFA, 8'hFA, 8'h20, 8'h21, 8'h21, 8'h61, 8'h21, 8'h01, 8'hB7, 8'hFF, 8'hBB, 8'h9A, 8'h97, 8'h01, 8'h01, 8'h61, 8'h21, 8'h21, 8'h62, 8'h22, 8'h62, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h61, 8'h21, 8'h21, 8'h21, 8'h20, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h01, 8'h01, 8'h01, 8'h00, 8'h01, 8'h01, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h62, 8'h21, 8'h62, 8'h61, 8'h61, 8'h22}, 
{8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h20, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h65, 8'h22}, 
{8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h62, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h22, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h62, 8'h62, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h21, 8'h22, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h61, 8'h20, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h20, 8'h21, 8'h21, 8'h61, 8'h22, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h22}, 
{8'h22, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h81, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h22, 8'h22, 8'h62, 8'h22, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h20, 8'h20, 8'h8D, 8'h20, 8'h20, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h20, 8'hFB, 8'h20, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'hBB, 8'h00, 8'h01, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h22}, 
{8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h81, 8'hC5, 8'hC5, 8'hA5, 8'hA5, 8'h60, 8'h61, 8'h61, 8'h61, 8'h61, 8'h22, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h22, 8'h62, 8'h22, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h60, 8'h8D, 8'h85, 8'hAD, 8'h20, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h20, 8'h20, 8'hFA, 8'hFA, 8'hFA, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h25, 8'h00, 8'hBB, 8'hBA, 8'hBB, 8'h01, 8'h01, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h80, 8'hC5, 8'hC5, 8'hC4, 8'hC4, 8'hC4, 8'hC5, 8'h60, 8'h60, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h22, 8'h21, 8'h22, 8'h22, 8'h21, 8'h01, 8'h01, 8'h26, 8'h01, 8'h22, 8'h21, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h22, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h20, 8'h85, 8'h60, 8'h60, 8'hFB, 8'hAD, 8'h20, 8'h21, 8'h21, 8'h61, 8'h21, 8'h20, 8'hFA, 8'h00, 8'h00, 8'hFF, 8'hFA, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'hBB, 8'h04, 8'h00, 8'hFF, 8'hBB, 8'h01, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h65, 8'h22}, 
{8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h81, 8'hC5, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hA5, 8'h60, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'hFF, 8'h85, 8'hA5, 8'hA5, 8'h21, 8'h01, 8'h21, 8'h21, 8'h22, 8'h01, 8'h05, 8'h05, 8'h0E, 8'h9B, 8'h9B, 8'hBB, 8'h01, 8'h21, 8'h22, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h62, 8'h21, 8'h61, 8'h61, 8'h20, 8'h8D, 8'hAD, 8'hAD, 8'h20, 8'h64, 8'h85, 8'h20, 8'h21, 8'h61, 8'h20, 8'h00, 8'hFA, 8'hFF, 8'hFA, 8'h00, 8'h00, 8'hFB, 8'h00, 8'h21, 8'h21, 8'h01, 8'h00, 8'hBB, 8'hBA, 8'hBA, 8'h00, 8'h00, 8'hBB, 8'h01, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h62, 8'h62, 8'h22, 8'h62, 8'h21, 8'h22}, 
{8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hCC, 8'hFA, 8'hC4, 8'hA4, 8'hA5, 8'h60, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'hFF, 8'hAD, 8'h85, 8'hAD, 8'h65, 8'h01, 8'h01, 8'h01, 8'h05, 8'h05, 8'h9B, 8'h7B, 8'h7B, 8'h9F, 8'h9B, 8'hBB, 8'h01, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h22, 8'h22, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h20, 8'h8D, 8'h20, 8'h20, 8'hFF, 8'hAD, 8'h20, 8'h20, 8'h20, 8'h21, 8'h21, 8'h00, 8'hFB, 8'h20, 8'h00, 8'hFF, 8'hFA, 8'h00, 8'h00, 8'h20, 8'h21, 8'h21, 8'h01, 8'hB7, 8'h04, 8'h04, 8'hFF, 8'hBA, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h22, 8'h22, 8'h62, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'hA5, 8'hC4, 8'hC4, 8'h60, 8'h60, 8'h60, 8'hA4, 8'hA4, 8'hC4, 8'hA5, 8'h60, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h21, 8'h61, 8'h20, 8'h61, 8'h20, 8'h20, 8'h00, 8'h05, 8'h76, 8'h9F, 8'h9F, 8'h7B, 8'h7F, 8'h3F, 8'h3F, 8'h3F, 8'h3B, 8'h05, 8'h05, 8'h21, 8'h21, 8'h20, 8'h61, 8'h61, 8'h81, 8'h81, 8'h61, 8'h61, 8'h61, 8'h22, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hAD, 8'h20, 8'h20, 8'h8D, 8'h20, 8'h20, 8'h21, 8'h61, 8'h21, 8'h20, 8'hFF, 8'hFA, 8'h00, 8'h00, 8'hFB, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h01, 8'hFF, 8'hBB, 8'h00, 8'h04, 8'hB6, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h21, 8'h21, 8'h65, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h60, 8'h60, 8'hC4, 8'hC4, 8'h60, 8'h60, 8'h60, 8'h60, 8'hC4, 8'hA4, 8'h60, 8'h60, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h20, 8'h20, 8'h00, 8'h00, 8'h04, 8'h04, 8'h76, 8'h9F, 8'h7A, 8'h3F, 8'h3F, 8'h3F, 8'h1F, 8'h1F, 8'h3F, 8'h3F, 8'h05, 8'h05, 8'hFF, 8'hFF, 8'h20, 8'h85, 8'hA5, 8'hA5, 8'hA5, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h20, 8'hFF, 8'h8D, 8'h00, 8'h20, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'hFF, 8'hFA, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h00, 8'hFF, 8'hBA, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h60, 8'hC4, 8'hC4, 8'hC4, 8'hA4, 8'hAC, 8'hFE, 8'hCC, 8'hA4, 8'h60, 8'h60, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'h60, 8'h60, 8'h20, 8'h00, 8'h00, 8'h00, 8'h9B, 8'h9A, 8'hBF, 8'hBF, 8'hBF, 8'hBF, 8'h9F, 8'h3F, 8'h1F, 8'h1F, 8'h1F, 8'h3F, 8'h7B, 8'hFF, 8'hFF, 8'hFF, 8'h20, 8'h85, 8'hAD, 8'hA5, 8'hAD, 8'h85, 8'h61, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h20, 8'h20, 8'h65, 8'h20, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'hDA, 8'h00, 8'h00, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h01, 8'h00, 8'hB6, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h22}, 
{8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h60, 8'h60, 8'hC4, 8'hC4, 8'hA4, 8'hAC, 8'h84, 8'hFF, 8'hA4, 8'hCD, 8'h20, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'hFF, 8'hA5, 8'hA5, 8'hA5, 8'h85, 8'h20, 8'h00, 8'h00, 8'h00, 8'h7A, 8'h9F, 8'h7A, 8'h7F, 8'hBF, 8'h7F, 8'h3A, 8'h3F, 8'h3F, 8'h1F, 8'h3F, 8'h7F, 8'h3A, 8'h04, 8'h00, 8'h00, 8'h00, 8'h20, 8'h60, 8'h60, 8'h60, 8'h60, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h62, 8'h22, 8'h62, 8'h21, 8'h21, 8'h21, 8'h20, 8'h20, 8'h00, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h00, 8'h20, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h01, 8'h01, 8'h00, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h22, 8'h62, 8'h22, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h22}, 
{8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h80, 8'hC4, 8'hC4, 8'h60, 8'h60, 8'h60, 8'hFF, 8'hAD, 8'h60, 8'h60, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'hFF, 8'hAD, 8'hA5, 8'hA5, 8'hAD, 8'h85, 8'h20, 8'h00, 8'h04, 8'h9F, 8'h7B, 8'h7F, 8'h9F, 8'h9F, 8'h9F, 8'h7F, 8'h3E, 8'h3F, 8'h3F, 8'h3F, 8'h3A, 8'hBF, 8'hDF, 8'hFF, 8'hFF, 8'h20, 8'h84, 8'hAD, 8'hAD, 8'hAD, 8'h85, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h00, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h62, 8'h21, 8'h62, 8'h21, 8'h65, 8'h21, 8'h22}, 
{8'h22, 8'h22, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hCD, 8'h80, 8'h60, 8'h60, 8'h20, 8'h60, 8'hAD, 8'hA5, 8'h60, 8'h60, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h20, 8'h60, 8'h60, 8'h85, 8'hAD, 8'h65, 8'h00, 8'h96, 8'h9B, 8'h7A, 8'hBF, 8'h9F, 8'h3A, 8'h9F, 8'h7F, 8'h7F, 8'h7F, 8'h7F, 8'h7A, 8'h0D, 8'hBF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h22, 8'h22, 8'h21, 8'h62, 8'h22, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h22}, 
{8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h81, 8'hC5, 8'hC4, 8'hC4, 8'hEC, 8'hC4, 8'hC4, 8'hCC, 8'hFA, 8'hCD, 8'hA5, 8'h81, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h60, 8'h20, 8'h20, 8'h00, 8'h01, 8'h00, 8'h05, 8'h9A, 8'h9B, 8'hDF, 8'hBF, 8'h0D, 8'h7A, 8'h9A, 8'h05, 8'h00, 8'h00, 8'h01, 8'h00, 8'h00, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h21, 8'h61, 8'h21, 8'h62, 8'h22, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h62, 8'h21, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h22}, 
{8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h81, 8'hC5, 8'hC4, 8'hC4, 8'hC4, 8'hC4, 8'hCC, 8'hA4, 8'hCC, 8'hA4, 8'hA5, 8'h60, 8'h61, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h01, 8'h01, 8'h00, 8'h00, 8'h01, 8'h97, 8'hBB, 8'h96, 8'h01, 8'h01, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h62, 8'h22, 8'h62, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h62, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h22, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hA4, 8'hCC, 8'hC4, 8'hC4, 8'hA4, 8'hCC, 8'hA4, 8'hCD, 8'hC5, 8'h60, 8'h61, 8'h21, 8'h21, 8'h62, 8'h62, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h01, 8'h21, 8'h21, 8'h01, 8'h26, 8'h01, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h62, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h61, 8'h21, 8'h62, 8'h21, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h62, 8'h21, 8'h61, 8'h61, 8'h61, 8'hA5, 8'hA5, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'hA5, 8'hA5, 8'h61, 8'h61, 8'h61, 8'h62, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h61, 8'h62, 8'h62, 8'h22, 8'h62, 8'h21, 8'h62, 8'h22, 8'h21, 8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'hFB, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h61, 8'h22}, 
{8'h62, 8'h62, 8'h22, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h22, 8'h22, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h20, 8'hFB, 8'hFB, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h21, 8'h22}, 
{8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h22, 8'h22, 8'h22, 8'h61, 8'h61, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h20, 8'hFA, 8'h20, 8'h20, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h21, 8'h61, 8'h21, 8'h65, 8'hFF, 8'h22}, 
{8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h21, 8'h61, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h20, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hD6, 8'h20, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h61, 8'h61, 8'hFF, 8'hFF, 8'h22}, 
{8'h61, 8'h61, 8'h21, 8'h21, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h61, 8'h61, 8'h62, 8'h62, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h21, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h21, 8'h61, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFF, 8'h00, 8'h21, 8'h61, 8'h21, 8'h21, 8'h61, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'h20, 8'h22}, 
{8'h22, 8'h21, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'h00, 8'h00, 8'h61, 8'h21, 8'h62, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h21, 8'h61, 8'hFF, 8'h21, 8'h22}, 
{8'h22, 8'h22, 8'h21, 8'h21, 8'h22, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h21, 8'h22, 8'h22, 8'h21, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h21, 8'h22, 8'h22, 8'h22, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h61, 8'h62, 8'h21, 8'h62, 8'h21, 8'h21, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hDA, 8'h00, 8'h00, 8'h20, 8'h21, 8'h21, 8'h62, 8'h22, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'hFF, 8'hFF, 8'h22}, 
{8'h22, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h22, 8'h61, 8'h61, 8'h62, 8'h62, 8'h21, 8'h21, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h22, 8'h62, 8'h61, 8'h61, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'h21, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFA, 8'h00, 8'h21, 8'h61, 8'h21, 8'h62, 8'h62, 8'h62, 8'h21, 8'h21, 8'h62, 8'h21, 8'h66, 8'hFB, 8'h22}, 
{8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h21, 8'h21, 8'h61, 8'h62, 8'h22, 8'h21, 8'h21, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h62, 8'h22, 8'h22, 8'h22, 8'h21, 8'h61, 8'h61, 8'h61, 8'h22, 8'h22, 8'h22, 8'h22, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h61, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h62, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h00, 8'h00, 8'hFF, 8'hFF, 8'h21, 8'h21, 8'h21, 8'h61, 8'h62, 8'h62, 8'h22, 8'h22, 8'h62, 8'h21, 8'h21, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h21, 8'h61, 8'h21, 8'h61, 8'h21, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'hFA, 8'hFA, 8'h00, 8'h21, 8'h21, 8'h62, 8'h21, 8'h21, 8'h61, 8'h21, 8'h62, 8'h21, 8'h61, 8'h21, 8'h61, 8'h22}, 
};

localparam  int BG_NUMBER_OF_Y_BITS = 1;  // 2^1 = 2 
localparam  int BG_NUMBER_OF_X_BITS = 8;  // 2^8 = 256 
localparam  int BG_HEIGHT_Y = 1 <<  BG_NUMBER_OF_Y_BITS ;
localparam  int BG_WIDTH_X = 1 <<  BG_NUMBER_OF_X_BITS;
localparam  int BG_HEIGHT_Y_DIVIDER = BG_NUMBER_OF_Y_BITS - 2; //how many pixel bits are in every collision pixel
localparam  int BG_WIDTH_X_DIVIDER =  BG_NUMBER_OF_X_BITS - 2;
//logic [0:BG_HEIGHT_Y-1] [0:BG_WIDTH_X-1] [7:0] background = {
//	{8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92},
//	{8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h15, 8'h15, 8'h15, 8'h15, 8'h15, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92, 8'h92},
//};
logic [0:31][0:127][7:0]  background = {
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h0c,8'h0c,8'h10,8'h34,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h30,8'h04,8'h04,8'h04,8'h04,8'h04,8'h2c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h74,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h0c,8'h04,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h78,8'h78,8'h78,8'h0c,8'h00,8'h04,8'h04,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h0c,8'h04,8'h04,8'h2c,8'h04,8'h0c,8'h04,8'h04,8'h00,8'h00,8'h78,8'h34,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h04,8'h30,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h0c,8'h00,8'h00,8'h0c,8'h00,8'h74,8'h30,8'h00,8'h00,8'h00,8'h10,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h74,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hbb,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h10,8'h0c,8'h99,8'h0c,8'h34,8'h0c,8'h78,8'h10,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h0c,8'hbe,8'h78,8'h79,8'h0c,8'h78,8'h04,8'h00,8'h00,8'h04,8'h74,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h9d,8'h9a,8'h2d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h99,8'h0c,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h7c,8'h00,8'h04,8'h30,8'h00,8'h00,8'h04,8'h30,8'h00,8'h04,8'h0c,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h10,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h04,8'h04,8'hbe,8'h00,8'h04,8'h04,8'h00,8'h00,8'h79,8'h38,8'h78,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h74,8'h78,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h30,8'h34,8'h00,8'h30,8'h04,8'h0c,8'h00,8'h30,8'h10,8'h78,8'h78,8'h78,8'h04,8'h2c,8'h04,8'h0c,8'h00,8'h78,8'h34,8'h10,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h2d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h0c,8'h04,8'h34,8'h0c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hbe,8'h9a,8'h04,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hbe,8'h04,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h04,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hbb,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h10,8'h30,8'h78,8'h78,8'h78,8'h34,8'h30,8'h78,8'h78,8'h30,8'h34,8'h78,8'h30,8'h74,8'h78,8'h78,8'h0c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h34,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h30,8'h34,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h2c,8'h2d,8'h00,8'h00,8'h2c,8'h78,8'h74,8'h2d,8'h00,8'h00,8'h04,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h74,8'h30,8'h30,8'h0c,8'h34,8'h78,8'h78,8'h70,8'h75,8'h00,8'h74,8'h38,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hbe,8'h9a,8'h24,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h9e,8'h04,8'h30,8'h78,8'h78,8'h78,8'h78,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h74,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h74,8'h74,8'h78,8'h78,8'h34,8'h38,8'h78,8'h74,8'h78,8'h78,8'h78,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h79,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h10,8'h30,8'h78,8'h78,8'h78,8'h78,8'h71,8'h2c,8'h00,8'h00,8'h74,8'h78,8'h75,8'h31,8'h04,8'h00,8'h0c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h00,8'h2c,8'h74,8'h0c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h71,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h0c,8'h31,8'h04,8'h00,8'h04,8'h78,8'h74,8'h2c,8'h04,8'h00,8'h04,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h04,8'h34,8'h30,8'h04,8'h00,8'h78,8'h74,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h79,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h78,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hbf,8'hba,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h34,8'h74,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h9d,8'h9a,8'h2d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h99,8'h0c,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h0c,8'h04,8'h04,8'h04,8'h04,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h10,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h04,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h34,8'h78,8'h78,8'h78,8'h34,8'h00,8'h30,8'h34,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h38,8'h04,8'h04,8'h04,8'h9a,8'h00,8'h04,8'h00,8'h00,8'h00,8'h0c,8'h78,8'h78,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h70,8'h04,8'h78,8'h78,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h04,8'h04,8'h00,8'h0c,8'h04,8'h78,8'h10,8'h00,8'h00,8'h04,8'h34,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hdf,8'h96,8'h00,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hdf,8'h00,8'h30,8'h78,8'h78,8'h78,8'h78,8'h0c,8'h0c,8'h9a,8'h0c,8'h0c,8'h0c,8'h34,8'h30,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h9e,8'h9a,8'h24,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h9e,8'h04,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h74,8'h75,8'h78,8'h0c,8'h74,8'h74,8'h0c,8'h04,8'h00,8'h04,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h74,8'h00,8'h30,8'h04,8'h04,8'h04,8'h0c,8'h04,8'h00,8'h04,8'h30,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h30,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h00,8'h2c,8'h70,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h78,8'h78,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h2c,8'h30,8'h78},
	{8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hba,8'h6d,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'h78,8'h10,8'h30,8'h78,8'h78,8'h78,8'h78,8'h78,8'h38,8'h0c,8'h30,8'h00,8'h74,8'h04,8'h2c,8'h00,8'h79,8'h0c,8'h78,8'h78,8'h78,8'h00,8'h00,8'h00,8'h00,8'h04,8'h30,8'h34,8'h04,8'h78,8'h78,8'h78},
	{8'h38,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h38,8'h38,8'h38,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78,8'hbe,8'h96,8'h04,8'h00,8'h2d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hdf,8'hbe,8'h04,8'h30,8'h38,8'h38,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h10,8'h04,8'h04,8'h04,8'h0c,8'h78,8'h78,8'h78,8'h78,8'h78,8'h10,8'h78,8'h10,8'h78,8'h10,8'h78,8'h78,8'h78,8'h78,8'h78,8'h78}};
int y_pos=0;


always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
			RGBout <= 1'b0;
	end
	
	else begin
		if(sprite_number==11'b0) begin
			RGBout <= object_colors[(requested_x-x_offset)/2][(requested_y-y_offset)/2];
		end
		// death_0
		else if(sprite_number==99) begin
			RGBout <= object_colors[32+(requested_x-x_offset)/2][(requested_y-y_offset)/2];
		end
		else if(sprite_number==100) begin
			RGBout <= object_colors[64+(requested_x-x_offset)/2][(requested_y-y_offset)/2];
		end
		else if(sprite_number==101) begin
			RGBout <= object_colors[96+(requested_x-x_offset)/2][(requested_y-y_offset)/2];
		end
		// death_1
		else if(sprite_number==102) begin
			RGBout <= object_colors[64-(requested_x+x_offset)/2][(requested_y-y_offset)/2];
		end
		else if(sprite_number==103) begin
			RGBout <= object_colors[96-(requested_x+x_offset)/2][(requested_y-y_offset)/2];
		end
		else if(sprite_number==104) begin
			RGBout <= object_colors[128-(requested_x+x_offset)/2][(requested_y-y_offset)/2];
		end

		else if(sprite_number==11'b1) begin
			RGBout <= object_colors[18+((requested_x-x_offset)/2)][57+((requested_y-y_offset)/2)];
		end
		else if(sprite_number==11'b11111) begin
			if((requested_x-x_offset)/4 < 128) begin
				RGBout <= background[((requested_y+y_offset)/4)%32][(requested_x-x_offset)/4];
			end
			else begin
				RGBout<= 8'b1111_1111;
			end
		end
		else begin
			RGBout <= 8'b1111_1111;
		end
	end
end

endmodule
