
const logic[0:15][0:15][7:0] ai_car_yellow = {
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'hf8,8'hff,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hf8,8'hff,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hff,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hff,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hff,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hff,8'h00,8'h00,8'h00,8'hf8,8'hf8,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h91,8'h00,8'h00,8'h00,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'hf8,8'hf8,8'hf8,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'hf8,8'hf8,8'hf8,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'hf8,8'hf8,8'hf8,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'hf8,8'hf8,8'hf8,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hf8,8'h00,8'h00,8'h00,8'hf8,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf8,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf8,8'h00,8'h00,8'h62,8'h62,8'h62}};

const logic[0:31][0:15][7:0] ai_truck = {
	{8'h62,8'h62,8'h62,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h00,8'h00,8'h00,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'hff,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h00,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h00,8'h00,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h1f,8'h00,8'h1f,8'h1f,8'h1f,8'h1f,8'h00,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h1f,8'hff,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h1f,8'hff,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h62},
	{8'h62,8'h62,8'h62,8'h00,8'h1f,8'h00,8'h00,8'h1f,8'h00,8'h00,8'h00,8'h62,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h62,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'h91,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00}};

logic[0:15][0:15][7:0] car_bonus_sprite = {
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h62,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hff,8'he4,8'he4,8'he4,8'he4,8'he4,8'hff,8'h00,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'hff,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hff,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'hff,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hff,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'hff,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'he4,8'hff,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'hff,8'he4,8'he4,8'h00,8'h00,8'h00,8'he4,8'he4,8'hff,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h62,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hff,8'h00,8'hf8,8'hf8,8'h1f,8'h00,8'hff,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hff,8'h00,8'hf8,8'hf8,8'h1f,8'h00,8'hff,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hff,8'hf8,8'hf8,8'hf8,8'h1f,8'h1f,8'hff,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'h00,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'hff,8'hf8,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'hff,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'hff,8'hf8,8'hf8,8'hf8,8'hf8,8'h1f,8'h1f,8'h1f,8'hff,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'hff,8'hf8,8'hf8,8'hf8,8'hf8,8'h1f,8'h1f,8'h1f,8'hff,8'h00,8'h00,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h62,8'h62,8'h62},
	{8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62,8'h62}};
