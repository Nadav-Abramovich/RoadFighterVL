reg hi;